C:\Users\Alan\source\repos\mididrums\schematics\mididrums.cir Transient Analysis
* Converted From Micro Cap Source file to PSPICE
*
.FUNC DPWR(D) {I(D)*V(D)}
.FUNC BPWR(Q) {IC(Q)*VCE(Q)+IB(Q)*VBE(Q)}
.FUNC FPWR(M) {ID(M)*VDS(M)}
.FUNC HOTD(D,MAX) {IF((V(D)*I(D)>MAX),1,0)}
.FUNC HOTB(Q,MAX) {IF((VCE(Q)*IC(Q)+IB(Q)*VBE(Q)>MAX),1,0)}
.FUNC HOTF(M,MAX) {IF((VDS(M)*ID(M)>MAX),1,0)}
.PARAM LOW3MIN={IMPORT(LOW3MIN.OUT,LOW3THRES)}
.PARAM HIGH3MAX={IMPORT(HIGH3MAX.OUT,HIGH3THRES)}
.PARAM LOWLVDS={IMPORT(LOWLVDS.OUT,LOWLIMIT)}
.PARAM HILVDS={IMPORT(HILVDS.OUT,HILIMIT)}
.PARAM LIMTLVDS={IMPORT(LIMTLVDS.OUT,LVDSLIMITS)}
.FUNC SKINAC(DCRES,RESISTIVITY,RELPERM,RADIUS) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHAC(RESISTIVITY,RELPERM))**2))*DCRES}
.FUNC SKINDEPTHAC(RESISTIVITY,RELPERM) {503.3*(SQRT(RESISTIVITY/(RELPERM*F)))}
.FUNC SKINTR(DCRES,RESISTIVITY,RELPERM,RADIUS,FREQ) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ))**2))*DCRES}
.FUNC SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ) {503.3*(SQRT(RESISTIVITY/(RELPERM*FREQ)))}
R1 1 2 50K
R4 4 0 100K
V1 1 0 DC 3.3 AC 0.5 0 
X1 3 4 0 4 1 $GENERIC
X2 0 3 2 POT PARAMS: POTSIZE=100K PERCENT=50 
*
*** From file C:\MC12\library\POT.MAC
.SUBCKT POT  PINA PINB PINC PARAMS: POTSIZE=10K PERCENT=50 
R1 PINB PINA {POTSIZE*PERCENT/100}
R2 PINC PINB {POTSIZE-R(R1)}
.ENDS POT
*
* OPAMP
* PINS:  1=NC+ 2=NC- 3=VEE 4=VO 5=VCC
.SUBCKT $GENERIC 1 2 3 4 5
RSUPPLUS 5 0 1
RSUPMIN  3 0 1
C1 6 0 0.000101859163578813
R1 6 0 125
G1 0 6 TABLE {V(1,2)} = (-0.3183098861837909,-0.1489190005519877)
+ (0.3183098861837909,0.1489190005519877)
C2 7 0 2.940454728735431e-010
R2 7 0 125
G2 0 7 6 0 0.4678428381140585
ROUT 4 0 125
GOUT 0 4 7 0 0.4678428381140585
RIN 1 2 1G
.ENDS $GENERIC
*
.OPTIONS ACCT LIST OPTS ABSTOL=1pA CHGTOL=.01pC DEFL=100u DEFW=100u DEFNRD=0
+ DEFNRS=0 DEFPD=0 DEFPS=0 DIGDRVF=2 DIGDRVZ=20K DIGERRDEFAULT=20 DIGERRLIMIT=0
+ DIGFREQ=10GHz DIGINITSTATE=0 DIGIOLVL=2 DIGMNTYMX=2 DIGMNTYSCALE=0.4 DIGOVRDRV=3
+ DIGTYMXSCALE=1.6 GMIN=1p ITL1=100 ITL2=50 ITL4=10 PIVREL=1m PIVTOL=.1p RELTOL=1m
+ TNOM=27 TRTOL=7 VNTOL=1u WIDTH=80
*
.LIB "C:\MC12\library\NOM.LIB"
*
.TEMP 27
*
.TRAN 0.0002 10m 0 
.PLOT TRAN v(1) v(2)
*
.PROBE
.END
;$SpiceType=PSPICE
